////////////////////////////////////////////////////////////////////////////////
//
// Lab 3 Memory Tester: Number to bitmap decoder
//
// This module converts a 4-bit input to a 80-dot (2 digit) bitmap representing
// the numbers ' 0' through '15'.
//
// Author: Yun Wu, Nathan Ickes
// Date: March 8, 2006
//
////////////////////////////////////////////////////////////////////////////////

module dots(clk, num, dots);
   input clk;
   input [3:0] num;
   output [79:0] dots;
   
   reg [79:0] dots;
   always @ (posedge clk)
     case (num)
       4'd15: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '15'
		       40'b00100111_01000101_01000101_01000101_00111001};
       4'd14: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '14'
		       40'b00011000_00010100_00010010_01111111_00010000};
       4'd13: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '13'
		       40'b00100010_01000001_01001001_01001001_00110110};
       4'd12: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '12'
		       40'b01100010_01010001_01001001_01001001_01000110};
       4'd11: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '11'
		       40'b00000000_01000010_01111111_01000000_00000000};
       4'd10: dots <= {40'b00000000_01000010_01111111_01000000_00000000, // '10'
		       40'b00111110_01010001_01001001_01000101_00111110};
       4'd09: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 9'
		       40'b00000110_01001001_01001001_00101001_00011110};
       4'd08: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 8'
		       40'b00110110_01001001_01001001_01001001_00110110};
       4'd07: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 7'
		       40'b00000001_01110001_00001001_00000101_00000011};
       4'd06: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 6'
		       40'b00111100_01001010_01001001_01001001_00110000};
       4'd05: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 5'
		       40'b00100111_01000101_01000101_01000101_00111001};
       4'd04: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 4'
		       40'b00011000_00010100_00010010_01111111_00010000};
       4'd03: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 3'
		       40'b00100010_01000001_01001001_01001001_00110110};
       4'd02: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 2'
		       40'b01100010_01010001_01001001_01001001_01000110};
       4'd01: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 1'
		       40'b00000000_01000010_01111111_01000000_00000000};
       4'd00: dots <= {40'b00000000_00000000_00000000_00000000_00000000, // ' 0'
		       40'b00111110_01010001_01001001_01000101_00111110};
       // No default case, becase every case is already accounted for.
     endcase
   
endmodule
